# Swedish
# Day names
S�n
M�n
Tis
Ons
Tor
Fre
L�r
# Months
Jan
Feb
Mar
Apr
Maj
Jun
Jul
Aug
Sep
Okt
Nov
Dec
# Additional labels
L�ge
GMT tid
Solst�nd
Nationell tid
Dagens l�ngd
Soluppg�ng
Solnedg�ng
#
sekunden
minut
timme
dag
dagar
#
Klicka p� en stad
Klicka p� en plats
Klicka p� tv� platser
Klick tv� g�nger eller sl� � f�r � ' "
#
Tastatur
Tastatur/Mus kontroll
Escape
Escape meny
Unknown key binding !!
Synchro
Tids-variabel =
Global tid variabel =
#
City name
Timezone
Latitude
Longitude
Size
Warning: %s, lat = %s lon = %s%salready in list of cities !!
Overriding previous entry for %s
#
Option
Activating selected option...
Option incorrect or not available at runtime !!
Options: strike <Ctrl><Space> for blank space within an item
(once)
(periodically, period %d seconds)
(with starry sky)
(blank root window)
with the following rather long list of options:
Starting from **, options are runtime configurable.
Calculating new image...
Sunclock har ett antal funktioner som kan �tkommas genom mus-klick eller tastaturet:
# General help
Visa hj�lp och alternativ (H eller mus-klick knapp 1)
Laddar karta Jord (F eller mus-klick knapp 2)
Zoom (Z eller mus-klick knapp 3)
Parameters of Urban locations
Option command window
Anv�nd koordinat mode
Anv�nd solst�nd mode
Anv�nd distans mode
Anv�nd timme extension mode
Anv�nd nationell tidszon mode
�ndra tiden Fram�t
�ndra tiden Bak�t
Justera tidsvariabel
�terst�ll Global tid
Rita/Radera Natt
Rita/Radera S�n och M�ne
Rita/Radera meridianer
Rita/Radera breddgrader
Rita/Radera Tropik/Ekvator/Arktik cirklar
�ppnar ny kartf�nster
Slutar f�nster
Ikonifiera f�nster
F�rnya kartf�nster
Adjust window width to screen size
Back till f�reg�ende kartf�nster m�tt
V�xla tidszon och kartf�nster 
Aktivera kommando (-command option)
Avsluta program
# Zoom window help
Activate new zoom settings
Return to previous zoom settings
Cancel change in zoom settings
Set aspect by resizing main window
Cycle through zoom modes 0,1,2
Zoom in by factor 1.2
Zoom out by factor 1/1.2 = 0.833
Return to zoom factor = 1 (full map)
Center zoom area on selected city or location
Synchronize zoom operation
# Option window help
Activate the option
Erase the option command line
Synchronize windows or not
Copy map to root window
Erase map from root window
Start/stop animation
# Urban window help
Use degrees, minutes, seconds, or decimal degrees
Search/select city
Modify city parameters
Create new city location
Delete city
# End
